module main

fn moves(discs int, poles int) int {
}
