module main

pub enum Category {
	ones
	twos
	threes
	fours
	fives
	sixes
	fullHouse
	fourOfAKind
	littleStraight
	bigStraight
	choice
	yacht
}

fn score(dice []int, category Category) int {
}
