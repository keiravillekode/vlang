module main

fn test_yacht() {
	assert score([5, 5, 5, 5, 5], .yacht) == 50
}

fn test_not_yacht() {
	assert score([1, 3, 3, 2, 5], .yacht) == 0
}

fn test_ones() {
	assert score([1, 1, 1, 3, 5], .ones) == 3
}

fn test_ones_out_of_order() {
	assert score([3, 1, 1, 5, 1], .ones) == 3
}

fn test_no_ones() {
	assert score([4, 3, 6, 5, 5], .ones) == 0
}

fn test_twos() {
	assert score([2, 3, 4, 5, 6], .twos) == 2
}

fn test_fours() {
	assert score([1, 4, 1, 4, 1], .fours) == 8
}

fn test_yacht_counted_as_threes() {
	assert score([3, 3, 3, 3, 3], .threes) == 15
}

fn test_yacht_of_3s_counted_as_fives() {
	assert score([3, 3, 3, 3, 3], .fives) == 0
}

fn test_fives() {
	assert score([1, 5, 3, 5, 3], .fives) == 10
}

fn test_sixes() {
	assert score([2, 3, 4, 5, 6], .sixes) == 6
}

fn test_full_house_two_small_three_big() {
	assert score([2, 2, 4, 4, 4], .full_house) == 16
}

fn test_full_house_three_small_two_big() {
	assert score([5, 3, 3, 5, 3], .full_house) == 19
}

fn test_two_pair_is_not_a_full_house() {
	assert score([2, 2, 4, 4, 5], .full_house) == 0
}

fn test_four_of_a_kind_is_not_a_full_house() {
	assert score([1, 4, 4, 4, 4], .full_house) == 0
}

fn test_yacht_is_not_a_full_house() {
	assert score([2, 2, 2, 2, 2], .full_house) == 0
}

fn test_four_of_a_kind() {
	assert score([6, 6, 4, 6, 6], .four_of_a_kind) == 24
}

fn test_yacht_can_be_scored_as_four_of_a_kind() {
	assert score([3, 3, 3, 3, 3], .four_of_a_kind) == 12
}

fn test_full_house_is_not_four_of_a_kind() {
	assert score([3, 3, 3, 5, 5], .four_of_a_kind) == 0
}

fn test_little_straight() {
	assert score([3, 5, 4, 1, 2], .little_straight) == 30
}

fn test_little_straight_as_big_straight() {
	assert score([1, 2, 3, 4, 5], .big_straight) == 0
}

fn test_four_in_order_but_not_a_little_straight() {
	assert score([1, 1, 2, 3, 4], .little_straight) == 0
}

fn test_no_pairs_but_not_a_little_straight() {
	assert score([1, 2, 3, 4, 6], .little_straight) == 0
}

fn test_minimum_is_1_maximum_is_5_but_not_a_little_straight() {
	assert score([1, 1, 3, 4, 5], .little_straight) == 0
}

fn test_big_straight() {
	assert score([4, 6, 2, 5, 3], .big_straight) == 30
}

fn test_big_straight_as_little_straight() {
	assert score([6, 5, 4, 3, 2], .little_straight) == 0
}

fn test_no_pairs_but_not_a_big_straight() {
	assert score([6, 5, 4, 3, 1], .big_straight) == 0
}

fn test_choice() {
	assert score([3, 3, 5, 6, 6], .choice) == 23
}

fn test_yacht_as_choice() {
	assert score([2, 2, 2, 2, 2], .choice) == 10
}
